`timescale 1ns/1ps

module test_mtvec_value;
  reg clk = 0;
  reg reset_n = 0;
  wire [31:0] pc_out;
  wire [31:0] instr_out;
  integer cycle_count = 0;

  always #5 clk = ~clk;

  rv32i_core_pipelined #(
    .RESET_VECTOR(32'h00000000),
    .MEM_FILE("tests/riscv-compliance/rv32ui-p-add.hex")
  ) dut (
    .clk(clk),
    .reset_n(reset_n),
    .pc_out(pc_out),
    .instr_out(instr_out)
  );

  always @(posedge clk) begin
    if (reset_n) begin
      cycle_count = cycle_count + 1;

      // Monitor mtvec writes around cycle 40-42
      if (dut.idex_csr_we && dut.idex_csr_addr == 12'h305) begin
        $display("Cycle %0d: Writing mtvec with value 0x%h at PC=%h",
                 cycle_count, dut.idex_csr_wdata, dut.idex_pc);
      end

      if (cycle_count >= 38 && cycle_count <= 44) begin
        $display("Cycle %0d: PC=%h mtvec=%h",
                 cycle_count, pc_out, dut.trap_vector);
      end

      if (cycle_count >= 46) $finish;
    end
  end

  initial begin
    #20 reset_n = 1;
  end
endmodule
