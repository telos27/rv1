// Floating-Point Compare Unit
// Implements FEQ.S/D, FLT.S/D, FLE.S/D instructions
// Pure combinational logic (1 cycle)
// Result written to integer register rd

`include "config/rv_config.vh"

module fp_compare #(
  parameter FLEN = `FLEN  // 32 for single-precision, 64 for double-precision
) (
  // Operands
  input  wire [FLEN-1:0]   operand_a,   // rs1
  input  wire [FLEN-1:0]   operand_b,   // rs2

  // Control (operation select)
  input  wire [1:0]        operation,   // 00: FEQ, 01: FLT, 10: FLE
  input  wire              fmt,          // 0: single-precision, 1: double-precision

  // Result (written to integer register)
  output reg  [31:0]       result,      // 0 or 1 (zero-extended to 32 bits)

  // Exception flags
  output reg               flag_nv      // Invalid operation (signaling NaN)
);

  // IEEE 754 format parameters
  localparam EXP_WIDTH = (FLEN == 32) ? 8 : 11;
  localparam MAN_WIDTH = (FLEN == 32) ? 23 : 52;

  // Extract components based on format
  // For FLEN=64 with single-precision (fmt=0): use bits [31:0] (NaN-boxed in [63:32])
  // For FLEN=64 with double-precision (fmt=1): use bits [63:0]
  // For FLEN=32: always single-precision
  wire sign_a;
  wire sign_b;
  wire [10:0] exp_a;  // Max exponent width (11 bits for double)
  wire [10:0] exp_b;
  wire [51:0] man_a;  // Max mantissa width (52 bits for double)
  wire [51:0] man_b;

  generate
    if (FLEN == 64) begin : g_flen64
      // For FLEN=64, support both single and double precision
      assign sign_a = fmt ? operand_a[63] : operand_a[31];
      assign sign_b = fmt ? operand_b[63] : operand_b[31];
      assign exp_a = fmt ? operand_a[62:52] : {3'b000, operand_a[30:23]};
      assign exp_b = fmt ? operand_b[62:52] : {3'b000, operand_b[30:23]};
      assign man_a = fmt ? operand_a[51:0] : {29'b0, operand_a[22:0]};
      assign man_b = fmt ? operand_b[51:0] : {29'b0, operand_b[22:0]};
    end else begin : g_flen32
      // For FLEN=32, only single-precision supported
      assign sign_a = operand_a[31];
      assign sign_b = operand_b[31];
      assign exp_a = {3'b000, operand_a[30:23]};
      assign exp_b = {3'b000, operand_b[30:23]};
      assign man_a = {29'b0, operand_a[22:0]};
      assign man_b = {29'b0, operand_b[22:0]};
    end
  endgenerate

  // Effective exponent/mantissa widths based on format
  wire [10:0] exp_all_ones = fmt ? 11'h7FF : 11'h0FF;  // All 1s for current format
  wire man_msb_a = fmt ? man_a[51] : man_a[22];         // MSB for NaN detection
  wire man_msb_b = fmt ? man_b[51] : man_b[22];

  // Detect special values
  wire is_nan_a = (exp_a == exp_all_ones) && (man_a != 0);
  wire is_nan_b = (exp_b == exp_all_ones) && (man_b != 0);
  wire is_snan_a = is_nan_a && !man_msb_a;  // Signaling NaN has MSB=0
  wire is_snan_b = is_nan_b && !man_msb_b;
  wire is_qnan_a = is_nan_a && man_msb_a;   // Quiet NaN has MSB=1
  wire is_qnan_b = is_nan_b && man_msb_b;

  // Check for zero (both +0 and -0) - exponent and mantissa both zero
  wire is_zero_a = (exp_a == 0) && (man_a == 0);
  wire is_zero_b = (exp_b == 0) && (man_b == 0);

  // Check for both zeros (+0 == -0 in IEEE 754)
  wire both_zero = is_zero_a && is_zero_b;

  // Floating-point comparison logic
  // Cannot use $signed() directly - FP format needs special handling!
  //
  // For FP comparison:
  // 1. If signs differ: negative < positive (unless both zero)
  // 2. If both positive: compare as unsigned (larger exp/mantissa = larger value)
  // 3. If both negative: compare as unsigned REVERSED (larger bit pattern = more negative = smaller value)

  wire both_positive = !sign_a && !sign_b;
  wire both_negative = sign_a && sign_b;
  wire signs_differ = sign_a != sign_b;

  // For positive numbers or when comparing magnitudes
  // Compare exponent first, then mantissa
  wire mag_a_less_than_b = (exp_a < exp_b) || ((exp_a == exp_b) && (man_a < man_b));
  wire a_equal_b = (sign_a == sign_b) && (exp_a == exp_b) && (man_a == man_b);

  // True FP less-than comparison
  wire a_less_than_b = both_zero ? 1'b0 :  // +0 and -0 are equal, not less than
                       signs_differ ? sign_a :  // If signs differ, negative (sign_a=1) < positive (sign_a=0)
                       both_positive ? mag_a_less_than_b :  // Both positive: normal magnitude compare
                       both_negative ? !mag_a_less_than_b && !a_equal_b : 1'b0;  // Both negative: reverse compare

  always @(*) begin
    // Default: no exception
    flag_nv = 1'b0;
    result = 32'd0;

    // Handle NaN cases
    if (is_nan_a || is_nan_b) begin
      case (operation)
        2'b00: begin  // FEQ
          // FEQ returns 0 for any NaN, no exception for quiet NaN
          result = 32'd0;
          flag_nv = is_snan_a || is_snan_b;  // Signal only if sNaN
        end
        2'b01, 2'b10: begin  // FLT, FLE
          // FLT/FLE return 0 for any NaN, always signal exception
          result = 32'd0;
          flag_nv = 1'b1;  // Always signal invalid for FLT/FLE with NaN
        end
        default: begin
          result = 32'd0;
          flag_nv = 1'b0;
        end
      endcase
    end
    // Handle normal comparison
    else begin
      case (operation)
        2'b00: begin  // FEQ: a == b
          // Special case: +0 == -0
          if (both_zero)
            result = 32'd1;
          else if (a_equal_b)
            result = 32'd1;
          else
            result = 32'd0;
        end
        2'b01: begin  // FLT: a < b
          // Special case: +0 and -0 are equal (not less than)
          if (both_zero)
            result = 32'd0;
          else if (a_less_than_b)
            result = 32'd1;
          else
            result = 32'd0;
        end
        2'b10: begin  // FLE: a <= b
          // Special case: +0 <= -0 is true
          if (both_zero)
            result = 32'd1;
          else if (a_less_than_b || a_equal_b)
            result = 32'd1;
          else
            result = 32'd0;
        end
        default: begin
          result = 32'd0;
        end
      endcase
    end
  end

endmodule
