`timescale 1ns/1ps

module test_csr_illegal;
  reg clk = 0;
  reg reset_n = 0;
  wire [31:0] pc_out;
  wire [31:0] instr_out;
  integer cycle_count = 0;

  always #5 clk = ~clk;

  rv32i_core_pipelined #(
    .RESET_VECTOR(32'h00000000),
    .MEM_FILE("tests/riscv-compliance/rv32ui-p-add.hex")
  ) dut (
    .clk(clk),
    .reset_n(reset_n),
    .pc_out(pc_out),
    .instr_out(instr_out)
  );

  always @(posedge clk) begin
    if (reset_n) begin
      cycle_count = cycle_count + 1;

      // Monitor CSR instruction and illegal_csr signal
      if (cycle_count >= 35 && cycle_count <= 40) begin
        $display("Cycle %0d: PC=%h", cycle_count, pc_out);
        $display("  idex_instr=%h idex_csr_addr=%h idex_csr_we=%b",
                 dut.idex_instruction, dut.idex_csr_addr, dut.idex_csr_we);
        $display("  ex_illegal_csr=%b idex_illegal_inst=%b idex_valid=%b",
                 dut.ex_illegal_csr, dut.idex_illegal_inst, dut.idex_valid);
        $display("  Combined illegal: (idex_illegal_inst | (ex_illegal_csr && idex_csr_we)) && idex_valid = %b",
                 (dut.idex_illegal_inst | (dut.ex_illegal_csr && dut.idex_csr_we)) && dut.idex_valid);
        $display("  exception=%b exception_code=%h", dut.exception, dut.exception_code);
        $display("");
      end

      if (cycle_count >= 42) $finish;
    end
  end

  initial begin
    #20 reset_n = 1;
  end
endmodule
